version https://git-lfs.github.com/spec/v1
oid sha256:732086076102ad5263bee2eeb3c9c97228366bfe03b73834bd25ea406dd0782d
size 3538
