version https://git-lfs.github.com/spec/v1
oid sha256:037d356e91bedc858e62abb1901474a2a9f284182af88e85c32db7e6eea1b165
size 13608
