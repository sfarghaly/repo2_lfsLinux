version https://git-lfs.github.com/spec/v1
oid sha256:76fddfa60686a42290308754fb6c4940264fd1f05c94216e0f64d7e47dc8938c
size 6191
