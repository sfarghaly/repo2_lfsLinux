version https://git-lfs.github.com/spec/v1
oid sha256:7dd1c6aa7eb14da70bb070cad087ad8dafc754b29e1c2ddc96e92e8ba4558c26
size 2285
