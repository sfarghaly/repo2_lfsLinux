version https://git-lfs.github.com/spec/v1
oid sha256:6ed625e48e7dc79a0ed5afc68c0ba28dcdd2920e5dd2d6f5b338cbfae9dacc60
size 831
