version https://git-lfs.github.com/spec/v1
oid sha256:3b9ba1a6b30848cd3baa0c69a13be961950b50d142c95bd1eabd7728ba7c203f
size 5794
