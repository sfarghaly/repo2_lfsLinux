version https://git-lfs.github.com/spec/v1
oid sha256:32e3d1f545b4b7dd9119aa557b4cda35662600b2d4612879eb6c7e9c0f778364
size 4150
