version https://git-lfs.github.com/spec/v1
oid sha256:d6b6211417fedeb5ee3f0459b225e6eb15fae82789a3e8c586199bea60cbf5d4
size 3924
