version https://git-lfs.github.com/spec/v1
oid sha256:7514d1f237a8ef8ac8fb5af2e4f2f61c7aea837b06e93266db65d3bede8b4e12
size 6594
