version https://git-lfs.github.com/spec/v1
oid sha256:f442e9126d3c59b0b2e0b5d77d91af9a366ec7fc2937c629fad5089df9c54b32
size 1250
