version https://git-lfs.github.com/spec/v1
oid sha256:2596f28a26d59cf58d45506aa26d2c4e77e34f6e3514c66150324d5187d18fad
size 5253
