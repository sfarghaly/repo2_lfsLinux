version https://git-lfs.github.com/spec/v1
oid sha256:f0e3e7b4a682e489a5fd5e78e0da9f4f75782652e70661b41e310fd536c37281
size 13437
