version https://git-lfs.github.com/spec/v1
oid sha256:97555c63c628b96ebe917da45179e9eec67d524b1432f8a2c567e4e66edd6671
size 1446
