version https://git-lfs.github.com/spec/v1
oid sha256:19e4156175a5b745b3fb8051cd65f9504af9a34ec9b43471db637e12068e5d51
size 11986
