version https://git-lfs.github.com/spec/v1
oid sha256:300bf6efc9e5a1a20139da5ad7f3a1a7b29e1e9022ec6182759dcbfae6208858
size 13714
