version https://git-lfs.github.com/spec/v1
oid sha256:52a1012a4890145ab889bd5f47b379b3b129c96799ef44a3b9e4d58f511ab3df
size 7502
