version https://git-lfs.github.com/spec/v1
oid sha256:deb1efab1ff30fd22ff92eea54867fba5f63b454509987f5dbad6dbc6575939c
size 6903
