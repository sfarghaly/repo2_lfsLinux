version https://git-lfs.github.com/spec/v1
oid sha256:03641f75c42a0522501bfc97234320d86c4b1eee5bedf953422a314c1e9b31e3
size 5131
