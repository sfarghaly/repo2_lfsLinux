version https://git-lfs.github.com/spec/v1
oid sha256:23e15eb6ceb8c971bbc50f96cf5c59e60f15b6dd514ff924ec2186494e194131
size 2607
