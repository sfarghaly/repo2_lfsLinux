version https://git-lfs.github.com/spec/v1
oid sha256:7c45abec5428e8ef79392f1af2883b2d62c8a63b33c17929439fba308ba55a61
size 46684
