version https://git-lfs.github.com/spec/v1
oid sha256:4366049df524e54ab5a506990e04bb1eabcd56d65afd5e647b1f333f71af2245
size 2761
