version https://git-lfs.github.com/spec/v1
oid sha256:9f2e1248a3e9ce7424106ffb7dbbf343e987419933b5f30818f178ba63d8ddf4
size 1972
