version https://git-lfs.github.com/spec/v1
oid sha256:af6171bea9f79c3f8ad702d3373b27f07c0b48d8f7df503242d2811c774c40a2
size 2672
