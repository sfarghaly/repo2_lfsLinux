version https://git-lfs.github.com/spec/v1
oid sha256:82c16942dbb2b95ef9af46741b759587cea652f063123a5c7d6ca7ae118eff99
size 6594
