version https://git-lfs.github.com/spec/v1
oid sha256:da64825e79f04dacdd1db8bb3226d34b2cc2881b5de801df5cb45243cc2d3555
size 14523
