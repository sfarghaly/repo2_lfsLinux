version https://git-lfs.github.com/spec/v1
oid sha256:1d6462816b17421e8edce061959037d48a6434f7ca29cbfdd97a8fc9ad4af946
size 1899
