version https://git-lfs.github.com/spec/v1
oid sha256:88210407f6feb24b27ca77a8d34469bef1b7cbedc7ff4dd16eb831c2d09e689a
size 16074
