version https://git-lfs.github.com/spec/v1
oid sha256:984ab33826e2146c244b03c9bdf66941c6bac8deef4ec381a9a17577cdb2d8cd
size 1665
