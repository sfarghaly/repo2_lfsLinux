version https://git-lfs.github.com/spec/v1
oid sha256:d926ff69ad082bddbdbf2cc3061e59e9299e85afda4d032d57aaf87b3ba818a8
size 73552
