version https://git-lfs.github.com/spec/v1
oid sha256:a94a7cba81b6f24f3078616b359071ee38efead54c0824792db9372d99bc3937
size 3361
