version https://git-lfs.github.com/spec/v1
oid sha256:7fb5b42a4cfcc5d82206a3cc8da9b8ca0810476a12fcf756b0f9d6d16c6ca829
size 8492
