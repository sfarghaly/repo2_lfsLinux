version https://git-lfs.github.com/spec/v1
oid sha256:54ba53a4bf7bd2d175037c9aa11135f45502ea062f821bce09aa8f053ff5d452
size 4178
