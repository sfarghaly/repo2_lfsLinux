version https://git-lfs.github.com/spec/v1
oid sha256:f618f75eef1d7adc9d9da2bfe193fdf18522d82e477f9108514e5bac957126e5
size 2715
