version https://git-lfs.github.com/spec/v1
oid sha256:93967f30c5a83e93922b75315a4166ed663ada83c8dbb9f6ba48ec3f3ce75745
size 1542
