version https://git-lfs.github.com/spec/v1
oid sha256:8853a44dcdb359dbb149ec8abb39a39ae44e3466cdc372943f31399b40ba8a91
size 10536
