version https://git-lfs.github.com/spec/v1
oid sha256:63992048bd943593feaa82ca5da2bd56edc598a930c65dc9517d88767dc7c9b3
size 6806
