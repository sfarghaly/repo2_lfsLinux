version https://git-lfs.github.com/spec/v1
oid sha256:38a3d6df559ea698298cc00963ae74afb9d211da6a3a74e136abfb23d66ed1ec
size 3035
