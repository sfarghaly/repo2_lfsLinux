version https://git-lfs.github.com/spec/v1
oid sha256:ee21dbb1aaf5b0af8c8892dcb6649a67a8d9a6bb285631f39966783f029347d5
size 4530
