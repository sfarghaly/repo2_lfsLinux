version https://git-lfs.github.com/spec/v1
oid sha256:9109bd284f6494b04712753d738ec67e6966aa18572b4702425fcc510fdc7218
size 7981
