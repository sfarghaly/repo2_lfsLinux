version https://git-lfs.github.com/spec/v1
oid sha256:527d13be8ea504b8f508f7dc08015921c2b67de3c6b48bd7063354db756158c5
size 2375
