version https://git-lfs.github.com/spec/v1
oid sha256:2e91c5fa4dcbf4c6f42d9b3222c27611e8a47fc4b85925bb6cc5769b8246b68c
size 3838
