version https://git-lfs.github.com/spec/v1
oid sha256:b6551cf890c06db06c66ebcd346a9922884a6da00494ef8d0869e341f0d0f6aa
size 4538
