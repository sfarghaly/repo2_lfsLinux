version https://git-lfs.github.com/spec/v1
oid sha256:49fd813a9fed98e1ed025799878c0fca49690a309434d5dae2a590b33de3078d
size 2145
