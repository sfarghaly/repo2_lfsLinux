version https://git-lfs.github.com/spec/v1
oid sha256:1d683b6e6c2b2a6f3c070fd232c562a4dd29857caea0ba5d23762efac700bc27
size 1667
