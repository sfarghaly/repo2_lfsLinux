version https://git-lfs.github.com/spec/v1
oid sha256:66593cba6be6d02e9bdc39f5f8b1e04e8ac42281117079e8728e83651bd6579e
size 6708
