version https://git-lfs.github.com/spec/v1
oid sha256:668da5d299aed66b84d3c72599f28188dc78c5c5658d30fdc9ddc01d4e12dbe9
size 4754
