version https://git-lfs.github.com/spec/v1
oid sha256:b8bea9219d9d6f8873e1eb9ebc9a4d8563100cebc29c959234ebfef4cf6e91a4
size 2178
