version https://git-lfs.github.com/spec/v1
oid sha256:7b87fd274a0e9fc65cf336c5a478afff6182f25c5b70b2a0f57036e5b1898045
size 2140
