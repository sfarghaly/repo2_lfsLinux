version https://git-lfs.github.com/spec/v1
oid sha256:521ff5f8947a397d9780c0d91d11dcb3bd4e1ef288133e14397f4d87e5f3e9f7
size 4201
