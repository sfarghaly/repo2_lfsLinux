version https://git-lfs.github.com/spec/v1
oid sha256:d03e2f75225bc9877ca7c1a5966905c2d2af5088ddbdd39ebe5b516e3ed2033f
size 4093
