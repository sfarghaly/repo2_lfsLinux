version https://git-lfs.github.com/spec/v1
oid sha256:0eb18f4ee2e7544fb696c219fb0880953cecb0c12ec768a5de7ce2c1f71752a4
size 867
