version https://git-lfs.github.com/spec/v1
oid sha256:9b50aa0db7cfa3b819088b6de39d379c71d5656e44fc5ee1a9bf56c8ccbf7bba
size 1937
