version https://git-lfs.github.com/spec/v1
oid sha256:2ada3bebc41c2e0d48a24b24e5ffc36cd720bef3a92c174947d065e5f948ee02
size 4190
