version https://git-lfs.github.com/spec/v1
oid sha256:76ae62a9af98b568674b7fe6273652bb2970440961a75476d4221e26ca790bb2
size 3521
