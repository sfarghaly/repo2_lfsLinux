version https://git-lfs.github.com/spec/v1
oid sha256:0fbd34f1c738f7ae36418ae091d90581b5c7f161965bf0427e55ed81f73d88d8
size 8095
