version https://git-lfs.github.com/spec/v1
oid sha256:fa8401b7d303902936c45ea689c32f29d9134d6c9b81770852e055f94904a160
size 2758
