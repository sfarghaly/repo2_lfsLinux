version https://git-lfs.github.com/spec/v1
oid sha256:381bda20567a5d6f5ad829ebb63d3bf4415f217adbe0e184e56ab869a3822e31
size 6005
