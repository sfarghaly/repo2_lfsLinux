version https://git-lfs.github.com/spec/v1
oid sha256:0e06716a84f28b24f99901f5a957b04abc53115395cebe2ccc663e7031914580
size 3597
