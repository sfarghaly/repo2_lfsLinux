version https://git-lfs.github.com/spec/v1
oid sha256:ac1212f387f99d305f7396b955dc3d78e2ce85d94e5069b3c53132d907470fdc
size 1805
