version https://git-lfs.github.com/spec/v1
oid sha256:0037aa10bf6be5d8f8e42dc792c55ee9258b8f0c50c6f0e563ff2664888f1853
size 13608
