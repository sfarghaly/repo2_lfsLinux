version https://git-lfs.github.com/spec/v1
oid sha256:cc8e70ff7d7d81c5a60a25d78954ddbdc5d995b9418db35027c8f00210757fb7
size 2748
