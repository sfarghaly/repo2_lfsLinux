version https://git-lfs.github.com/spec/v1
oid sha256:0f51656efbd7c2e57720b75bb8b99d6d9414792f66dab027b351ccdf031253e9
size 8206
