version https://git-lfs.github.com/spec/v1
oid sha256:3befa982e479bea3508a885b2f273e35ea6fa209780541d63d4091411c671a51
size 2078
