version https://git-lfs.github.com/spec/v1
oid sha256:4ef00b9506e1799224370fea0500a92e802c06773e0a48733b37205e962e122f
size 15478
