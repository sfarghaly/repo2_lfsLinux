version https://git-lfs.github.com/spec/v1
oid sha256:fb18130ad979d7c3b6895a73cbec2e57e70b4314315473dd9e72bee619ac2dad
size 3521
