version https://git-lfs.github.com/spec/v1
oid sha256:9966ad8dbc8f017b00098ea788388564f4c6983a2668b4a791dba99abbc0c1f6
size 7981
