version https://git-lfs.github.com/spec/v1
oid sha256:b115a68ac1dbd84bf62ef71e1b10392fd2bac3d8dfa98be30568f26ea798f6e7
size 2672
