version https://git-lfs.github.com/spec/v1
oid sha256:545dfe437f420ae09ff03e9a1f1aa322f1a4b92e3b4b915bef99dc596b770d79
size 6708
