version https://git-lfs.github.com/spec/v1
oid sha256:48f11163b81a5628d59646e9bc1530eb8371f6ca47be98d2e3587fd118f6bab1
size 2667
