version https://git-lfs.github.com/spec/v1
oid sha256:6bbbae11d22f465119898de9b25f555d8b3ca21419d013407571a5e354ceeb95
size 5419
