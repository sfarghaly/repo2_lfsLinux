version https://git-lfs.github.com/spec/v1
oid sha256:8a3058b291af3a4147ca08d98f484769aee47e0f2c0cdbb0e59dfbd3e5e84137
size 2596
