version https://git-lfs.github.com/spec/v1
oid sha256:e6b23787a8735550e0761aababe833683a844d4104b3e9e92319527b52add209
size 7707
