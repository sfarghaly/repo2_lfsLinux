version https://git-lfs.github.com/spec/v1
oid sha256:db7c937690c72108d144a969c895c24dc1a2ed28ad3826ea95b3d55accae58cc
size 2084
