version https://git-lfs.github.com/spec/v1
oid sha256:ec180ca599d1c1128f3bef9cd949f6993d2fd7794fdafcca6b3c5f0fed9d34f3
size 3596
