version https://git-lfs.github.com/spec/v1
oid sha256:85aee8769e38f7eb575105820bde2c66ba4ff12f7758721b23ef0788880f6d84
size 2744
