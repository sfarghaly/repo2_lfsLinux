version https://git-lfs.github.com/spec/v1
oid sha256:a9b9ec53dc58988c940da8505a672a26d3be9e2520819497cc7afaa7b9894a68
size 1490
