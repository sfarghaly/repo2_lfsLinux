version https://git-lfs.github.com/spec/v1
oid sha256:e692f7efc57c70c3ba9729edf3b47c1072100386e41b590e795ff67b2634f96c
size 3780
