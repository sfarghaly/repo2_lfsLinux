version https://git-lfs.github.com/spec/v1
oid sha256:2f62c1ee128bca9a704695e75e16d4439b0392145dae9ad26b22a79d0ba37265
size 4093
