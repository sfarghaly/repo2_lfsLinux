version https://git-lfs.github.com/spec/v1
oid sha256:1d87eddd91592c67dddcfd3870846d2d6d621aeadae2f0937c7bed63874c94d3
size 1505
