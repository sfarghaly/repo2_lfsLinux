version https://git-lfs.github.com/spec/v1
oid sha256:01624a6ab0015d6da4ca5f3514d654dba84d99c7c340285f76546a79130baaac
size 4447
