version https://git-lfs.github.com/spec/v1
oid sha256:9378ab0522bad01bb28ce77e572416f18ad75db5c8703432fb6645f4a90057b5
size 1695
