version https://git-lfs.github.com/spec/v1
oid sha256:8d23702b42d924342793a0b83ed31256419b372dd7d50a612411f0e5c1539b8f
size 2254
