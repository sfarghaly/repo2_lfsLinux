version https://git-lfs.github.com/spec/v1
oid sha256:5ba45fbd0d2fa550e8b7ea8c133a4ddd344ebe3870f17edbc867bf00986c4634
size 5499
