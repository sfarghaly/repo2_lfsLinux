version https://git-lfs.github.com/spec/v1
oid sha256:0d333613e6c72632f653a5c554f2807036c35673e32f7b76d0bb161e1740217c
size 2140
