version https://git-lfs.github.com/spec/v1
oid sha256:71ce4a79b9886e4c3d9794b7f01fd0125dc465f8a7b392e9715b39428d725806
size 1988
