version https://git-lfs.github.com/spec/v1
oid sha256:707df10917dfc09504b2a88e73f779050bbe84dfafbdbf7c2b6cfbac419efe18
size 9776
