version https://git-lfs.github.com/spec/v1
oid sha256:0ba898e8b02da11c226d52e984713d9a9082c29878ffe6bc3c65e9f6b0ca67d4
size 1451
