version https://git-lfs.github.com/spec/v1
oid sha256:2227d5d53b108047a65760fd5cbed025513eedcc18a6767442072353d90f3352
size 2761
