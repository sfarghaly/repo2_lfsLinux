version https://git-lfs.github.com/spec/v1
oid sha256:25bf8af00b27299aeb7edf731a5e7712eb89cb043843ba5e6fcc8e681843119c
size 3356
