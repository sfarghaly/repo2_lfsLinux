version https://git-lfs.github.com/spec/v1
oid sha256:ec927e3606d60ab60bc0cbe428b8cbf14e2180cdfc7ae034a24012a7c5c5cc69
size 4819
