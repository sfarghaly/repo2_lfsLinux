version https://git-lfs.github.com/spec/v1
oid sha256:e3d9d578bd977b7890bf1da62ca932431a8dc7bec9a625fc8f10ce79f33c69c8
size 12578
