version https://git-lfs.github.com/spec/v1
oid sha256:4d1ea4801c8906edc7f659f53ca865405b0b23ccb3e5e1b3ee155b2c0339a15f
size 2827
