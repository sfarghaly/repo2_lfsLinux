version https://git-lfs.github.com/spec/v1
oid sha256:77641decd95973f2c0cd7dafd2474989c66be17f918a205c1feff53d800d72d2
size 1184
