version https://git-lfs.github.com/spec/v1
oid sha256:3dc63c4140194add46385f03360ca8cfe6f094cf6e14a4318166be96fe0f059e
size 27281
