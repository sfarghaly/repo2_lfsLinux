version https://git-lfs.github.com/spec/v1
oid sha256:b16b6b582e17d5a511b5b4832cfa1325b968e4d5f0ac56427c3abd4f1b5dd4e7
size 2084
