version https://git-lfs.github.com/spec/v1
oid sha256:87795c47a2fcb56ef653229c44708e953d6482f9ecf5eee0878885848212d1d1
size 12220
