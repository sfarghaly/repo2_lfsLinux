version https://git-lfs.github.com/spec/v1
oid sha256:9ae845e6d7b52f9192e7fb711e5bd8ddf350b8349479fb52c531c648dc51d90d
size 3328
