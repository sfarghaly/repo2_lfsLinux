version https://git-lfs.github.com/spec/v1
oid sha256:d5147551099b7ae90bce2d6864aa84e4c9619252df1c76b84a439a2e0132bc9c
size 6151
