version https://git-lfs.github.com/spec/v1
oid sha256:86c1d06628c06b9d2dc14d75681b9f8ba5c4f1cc04f678325ae083175a71d900
size 2375
