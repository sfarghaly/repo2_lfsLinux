version https://git-lfs.github.com/spec/v1
oid sha256:dd8c60f84508d03e353bd16991fba95249da7408fad673da1a4c4ad3c50aa77c
size 5981
