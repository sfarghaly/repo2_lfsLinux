version https://git-lfs.github.com/spec/v1
oid sha256:b2354be0687a76e542e6fc57c764a803c784015300067c00717c058b1f60f358
size 3227
